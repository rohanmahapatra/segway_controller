library verilog;
use verilog.vl_types.all;
entity ISOLOD4BWP is
    port(
        ISO             : in     vl_logic;
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end ISOLOD4BWP;
