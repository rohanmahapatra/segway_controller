library verilog;
use verilog.vl_types.all;
entity GBUFFD2BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end GBUFFD2BWP;
