library verilog;
use verilog.vl_types.all;
entity GDFQD1BWP is
    port(
        D               : in     vl_logic;
        CP              : in     vl_logic;
        Q               : out    vl_logic
    );
end GDFQD1BWP;
