library verilog;
use verilog.vl_types.all;
entity OD25DCAP32BWP is
end OD25DCAP32BWP;
