library verilog;
use verilog.vl_types.all;
entity DCAPX8BWP is
end DCAPX8BWP;
