library verilog;
use verilog.vl_types.all;
entity EDFCNQD2BWP is
    port(
        D               : in     vl_logic;
        E               : in     vl_logic;
        CP              : in     vl_logic;
        CDN             : in     vl_logic;
        Q               : out    vl_logic
    );
end EDFCNQD2BWP;
