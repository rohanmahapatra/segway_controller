library verilog;
use verilog.vl_types.all;
entity LVLLHD4BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end LVLLHD4BWP;
