library verilog;
use verilog.vl_types.all;
entity XOR2D1BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        Z               : out    vl_logic
    );
end XOR2D1BWP;
