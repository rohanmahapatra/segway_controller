library verilog;
use verilog.vl_types.all;
entity DFCNQD2BWP is
    port(
        D               : in     vl_logic;
        CP              : in     vl_logic;
        CDN             : in     vl_logic;
        Q               : out    vl_logic
    );
end DFCNQD2BWP;
