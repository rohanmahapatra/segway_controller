library verilog;
use verilog.vl_types.all;
entity DEL225D1BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DEL225D1BWP;
