library verilog;
use verilog.vl_types.all;
entity GFILL4BWP is
end GFILL4BWP;
