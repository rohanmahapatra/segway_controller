library verilog;
use verilog.vl_types.all;
entity LVLLHD8BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end LVLLHD8BWP;
