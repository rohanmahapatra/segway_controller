library verilog;
use verilog.vl_types.all;
entity ND3D4BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        ZN              : out    vl_logic
    );
end ND3D4BWP;
