library verilog;
use verilog.vl_types.all;
entity CKND20BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end CKND20BWP;
