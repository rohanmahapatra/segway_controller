library verilog;
use verilog.vl_types.all;
entity INR2XD1BWP is
    port(
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        ZN              : out    vl_logic
    );
end INR2XD1BWP;
