library verilog;
use verilog.vl_types.all;
entity BHDBWP is
    port(
        Z               : inout  vl_logic
    );
end BHDBWP;
