library verilog;
use verilog.vl_types.all;
entity CKBD24BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end CKBD24BWP;
