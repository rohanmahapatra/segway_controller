library verilog;
use verilog.vl_types.all;
entity INR4D4BWP is
    port(
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        ZN              : out    vl_logic
    );
end INR4D4BWP;
