library verilog;
use verilog.vl_types.all;
entity GFILL3BWP is
end GFILL3BWP;
