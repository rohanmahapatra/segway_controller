library verilog;
use verilog.vl_types.all;
entity DCAPBWP is
end DCAPBWP;
