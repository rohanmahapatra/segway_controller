library verilog;
use verilog.vl_types.all;
entity DEL1D1BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DEL1D1BWP;
