library verilog;
use verilog.vl_types.all;
entity BUFFD3BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end BUFFD3BWP;
