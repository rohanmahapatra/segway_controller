library verilog;
use verilog.vl_types.all;
entity GFILL10BWP is
end GFILL10BWP;
