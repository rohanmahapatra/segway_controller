library verilog;
use verilog.vl_types.all;
entity DCCKBD20BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DCCKBD20BWP;
