library verilog;
use verilog.vl_types.all;
entity DCCKND20BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end DCCKND20BWP;
