library verilog;
use verilog.vl_types.all;
entity DCCKBD8BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DCCKBD8BWP;
