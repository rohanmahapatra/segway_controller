library verilog;
use verilog.vl_types.all;
entity DEL500D1BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DEL500D1BWP;
