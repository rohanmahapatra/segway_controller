library verilog;
use verilog.vl_types.all;
entity DEL075D1BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DEL075D1BWP;
