library verilog;
use verilog.vl_types.all;
entity GTIEHBWP is
    port(
        Z               : out    vl_logic
    );
end GTIEHBWP;
