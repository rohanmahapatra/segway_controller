library verilog;
use verilog.vl_types.all;
entity GOR2D2BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        Z               : out    vl_logic
    );
end GOR2D2BWP;
