library verilog;
use verilog.vl_types.all;
entity LVLHLD8BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end LVLHLD8BWP;
