library verilog;
use verilog.vl_types.all;
entity INVD2BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end INVD2BWP;
