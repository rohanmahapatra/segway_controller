// to be filled 
