library verilog;
use verilog.vl_types.all;
entity GTIELBWP is
    port(
        ZN              : out    vl_logic
    );
end GTIELBWP;
