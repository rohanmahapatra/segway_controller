library verilog;
use verilog.vl_types.all;
entity DCAPX64BWP is
end DCAPX64BWP;
