library verilog;
use verilog.vl_types.all;
entity LVLHLD2BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end LVLHLD2BWP;
