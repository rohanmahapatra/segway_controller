library verilog;
use verilog.vl_types.all;
entity GINVD1BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end GINVD1BWP;
