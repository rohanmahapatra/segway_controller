library verilog;
use verilog.vl_types.all;
entity DFQD1BWP is
    port(
        D               : in     vl_logic;
        CP              : in     vl_logic;
        Q               : out    vl_logic
    );
end DFQD1BWP;
