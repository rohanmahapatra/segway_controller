library verilog;
use verilog.vl_types.all;
entity INVD24BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end INVD24BWP;
