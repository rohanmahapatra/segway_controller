library verilog;
use verilog.vl_types.all;
entity OD25DCAP64BWP is
end OD25DCAP64BWP;
