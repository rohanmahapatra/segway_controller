library verilog;
use verilog.vl_types.all;
entity OD25DCAP16BWP is
end OD25DCAP16BWP;
