library verilog;
use verilog.vl_types.all;
entity DCAP64BWP is
end DCAP64BWP;
