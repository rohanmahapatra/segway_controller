library verilog;
use verilog.vl_types.all;
entity OA221D4BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        C               : in     vl_logic;
        Z               : out    vl_logic
    );
end OA221D4BWP;
