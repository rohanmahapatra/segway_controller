library verilog;
use verilog.vl_types.all;
entity GINVD3BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end GINVD3BWP;
