library verilog;
use verilog.vl_types.all;
entity CKND16BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end CKND16BWP;
