library verilog;
use verilog.vl_types.all;
entity GDCAP4BWP is
end GDCAP4BWP;
