library verilog;
use verilog.vl_types.all;
entity INVD3BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end INVD3BWP;
