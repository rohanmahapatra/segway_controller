library verilog;
use verilog.vl_types.all;
entity DCAP32BWP is
end DCAP32BWP;
