library verilog;
use verilog.vl_types.all;
entity AO31D1BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        B               : in     vl_logic;
        Z               : out    vl_logic
    );
end AO31D1BWP;
