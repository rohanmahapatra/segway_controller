library verilog;
use verilog.vl_types.all;
entity XNR3D2BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        ZN              : out    vl_logic
    );
end XNR3D2BWP;
