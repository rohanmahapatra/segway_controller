library verilog;
use verilog.vl_types.all;
entity DCAPX32BWP is
end DCAPX32BWP;
