library verilog;
use verilog.vl_types.all;
entity OR4XD1BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        A4              : in     vl_logic;
        Z               : out    vl_logic
    );
end OR4XD1BWP;
