library verilog;
use verilog.vl_types.all;
entity OA211D0BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        Z               : out    vl_logic
    );
end OA211D0BWP;
