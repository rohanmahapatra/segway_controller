library verilog;
use verilog.vl_types.all;
entity OR2D0BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        Z               : out    vl_logic
    );
end OR2D0BWP;
