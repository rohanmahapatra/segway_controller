library verilog;
use verilog.vl_types.all;
entity CKND24BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end CKND24BWP;
