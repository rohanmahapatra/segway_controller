library verilog;
use verilog.vl_types.all;
entity CKBD3BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end CKBD3BWP;
