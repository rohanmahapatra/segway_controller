library verilog;
use verilog.vl_types.all;
entity DCAP8BWP is
end DCAP8BWP;
