library verilog;
use verilog.vl_types.all;
entity DCCKBD4BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DCCKBD4BWP;
