library verilog;
use verilog.vl_types.all;
entity LVLHLD1BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end LVLHLD1BWP;
