library verilog;
use verilog.vl_types.all;
entity CKND1BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end CKND1BWP;
