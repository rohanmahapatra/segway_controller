library verilog;
use verilog.vl_types.all;
entity GDCAP2BWP is
end GDCAP2BWP;
