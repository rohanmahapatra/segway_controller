library verilog;
use verilog.vl_types.all;
entity GDCAPBWP is
end GDCAPBWP;
