library verilog;
use verilog.vl_types.all;
entity LVLHLD4BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end LVLHLD4BWP;
