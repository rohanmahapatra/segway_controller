library verilog;
use verilog.vl_types.all;
entity AN2D1BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        Z               : out    vl_logic
    );
end AN2D1BWP;
