library verilog;
use verilog.vl_types.all;
entity DCAP4BWP is
end DCAP4BWP;
