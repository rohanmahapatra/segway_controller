library verilog;
use verilog.vl_types.all;
entity AOI21D1BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B               : in     vl_logic;
        ZN              : out    vl_logic
    );
end AOI21D1BWP;
