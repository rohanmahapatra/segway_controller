library verilog;
use verilog.vl_types.all;
entity GOAI21D1BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B               : in     vl_logic;
        ZN              : out    vl_logic
    );
end GOAI21D1BWP;
