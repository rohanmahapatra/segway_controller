library verilog;
use verilog.vl_types.all;
entity INVD1BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end INVD1BWP;
