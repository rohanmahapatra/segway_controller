library verilog;
use verilog.vl_types.all;
entity AOI211D4BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        ZN              : out    vl_logic
    );
end AOI211D4BWP;
