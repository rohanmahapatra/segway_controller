library verilog;
use verilog.vl_types.all;
entity DCCKND16BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end DCCKND16BWP;
