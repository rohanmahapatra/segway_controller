library verilog;
use verilog.vl_types.all;
entity ANTENNABWP is
    port(
        I               : in     vl_logic
    );
end ANTENNABWP;
