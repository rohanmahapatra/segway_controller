library verilog;
use verilog.vl_types.all;
entity GDCAP3BWP is
end GDCAP3BWP;
