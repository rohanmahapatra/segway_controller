library verilog;
use verilog.vl_types.all;
entity GFILL2BWP is
end GFILL2BWP;
