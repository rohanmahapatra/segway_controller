library verilog;
use verilog.vl_types.all;
entity DEL125D1BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DEL125D1BWP;
