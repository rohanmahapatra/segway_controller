library verilog;
use verilog.vl_types.all;
entity GBUFFD4BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end GBUFFD4BWP;
