library verilog;
use verilog.vl_types.all;
entity DFXQD1BWP is
    port(
        DA              : in     vl_logic;
        DB              : in     vl_logic;
        SA              : in     vl_logic;
        CP              : in     vl_logic;
        Q               : out    vl_logic
    );
end DFXQD1BWP;
