library verilog;
use verilog.vl_types.all;
entity TIEHBWP is
    port(
        Z               : out    vl_logic
    );
end TIEHBWP;
