library verilog;
use verilog.vl_types.all;
entity DCAPX4BWP is
end DCAPX4BWP;
