library verilog;
use verilog.vl_types.all;
entity DCAP16BWP is
end DCAP16BWP;
