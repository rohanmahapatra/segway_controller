library verilog;
use verilog.vl_types.all;
entity OA33D2BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        Z               : out    vl_logic
    );
end OA33D2BWP;
