library verilog;
use verilog.vl_types.all;
entity BUFFD1BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end BUFFD1BWP;
