library verilog;
use verilog.vl_types.all;
entity NR2D4BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        ZN              : out    vl_logic
    );
end NR2D4BWP;
