library verilog;
use verilog.vl_types.all;
entity tsmc_xbuf is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end tsmc_xbuf;
