library verilog;
use verilog.vl_types.all;
entity DCAPX16BWP is
end DCAPX16BWP;
