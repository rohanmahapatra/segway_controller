library verilog;
use verilog.vl_types.all;
entity TIELBWP is
    port(
        ZN              : out    vl_logic
    );
end TIELBWP;
