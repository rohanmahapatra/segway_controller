library verilog;
use verilog.vl_types.all;
entity GFILLBWP is
end GFILLBWP;
