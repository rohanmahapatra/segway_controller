library verilog;
use verilog.vl_types.all;
entity CKLNQD3BWP is
    port(
        TE              : in     vl_logic;
        E               : in     vl_logic;
        CP              : in     vl_logic;
        Q               : out    vl_logic
    );
end CKLNQD3BWP;
