library verilog;
use verilog.vl_types.all;
entity LHQD2BWP is
    port(
        D               : in     vl_logic;
        E               : in     vl_logic;
        Q               : out    vl_logic
    );
end LHQD2BWP;
