library verilog;
use verilog.vl_types.all;
entity MOAI22D1BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        ZN              : out    vl_logic
    );
end MOAI22D1BWP;
