library verilog;
use verilog.vl_types.all;
entity GBUFFD3BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end GBUFFD3BWP;
