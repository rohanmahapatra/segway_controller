library verilog;
use verilog.vl_types.all;
entity IOA21D4BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B               : in     vl_logic;
        ZN              : out    vl_logic
    );
end IOA21D4BWP;
