library verilog;
use verilog.vl_types.all;
entity DCCKBD16BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end DCCKBD16BWP;
