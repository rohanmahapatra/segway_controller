library verilog;
use verilog.vl_types.all;
entity BUFFD2BWP is
    port(
        I               : in     vl_logic;
        Z               : out    vl_logic
    );
end BUFFD2BWP;
