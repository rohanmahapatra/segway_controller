library verilog;
use verilog.vl_types.all;
entity AN4D8BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        A4              : in     vl_logic;
        Z               : out    vl_logic
    );
end AN4D8BWP;
