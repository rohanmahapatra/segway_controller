library verilog;
use verilog.vl_types.all;
entity MAOI222D2BWP is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        ZN              : out    vl_logic
    );
end MAOI222D2BWP;
