library verilog;
use verilog.vl_types.all;
entity INVD0BWP is
    port(
        I               : in     vl_logic;
        ZN              : out    vl_logic
    );
end INVD0BWP;
