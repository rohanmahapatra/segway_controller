library verilog;
use verilog.vl_types.all;
entity OAI221D0BWP is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        C               : in     vl_logic;
        ZN              : out    vl_logic
    );
end OAI221D0BWP;
