library verilog;
use verilog.vl_types.all;
entity GDCAP10BWP is
end GDCAP10BWP;
