library verilog;
use verilog.vl_types.all;
entity INR3D2BWP is
    port(
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        ZN              : out    vl_logic
    );
end INR3D2BWP;
